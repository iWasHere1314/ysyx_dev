`include "defines.v"
module ex2mem(
    
);
    
endmodule